module top(input logic clk, reset,
	   output logic [31:0] writedata, dataadr,
	   output logic memwrite);

logic [31:0] pc, instr, readdata;
logic sb;		//To choose whether L'B', L'W'

// instantiate processor and memories
mips mips(clk, reset, pc, instr, memwrite, sb, dataadr, writedata, readdata);

imem imem(pc[7:2], instr);

dmem dmem(clk, memwrite, sb, dataadr, writedata, readdata);
endmodule
